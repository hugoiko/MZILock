


module red_pitaya_top (
   // PS connections
   inout  wire  [54-1: 0] FIXED_IO_mio       ,
   inout  wire            FIXED_IO_ps_clk    ,
   inout  wire            FIXED_IO_ps_porb   ,
   inout  wire            FIXED_IO_ps_srstb  ,
   inout  wire            FIXED_IO_ddr_vrn   ,
   inout  wire            FIXED_IO_ddr_vrp   ,
   // DDR
   inout  wire  [15-1: 0] DDR_addr           ,
   inout  wire  [ 3-1: 0] DDR_ba             ,
   inout  wire            DDR_cas_n          ,
   inout  wire            DDR_ck_n           ,
   inout  wire            DDR_ck_p           ,
   inout  wire            DDR_cke            ,
   inout  wire            DDR_cs_n           ,
   inout  wire  [ 4-1: 0] DDR_dm             ,
   inout  wire  [32-1: 0] DDR_dq             ,
   inout  wire  [ 4-1: 0] DDR_dqs_n          ,
   inout  wire  [ 4-1: 0] DDR_dqs_p          ,
   inout  wire            DDR_odt            ,
   inout  wire            DDR_ras_n          ,
   inout  wire            DDR_reset_n        ,
   inout  wire            DDR_we_n           ,

   // Red Pitaya periphery
  
   // ADC
   input  wire  [16-1: 2] adc_dat_a_i        ,  // ADC CH1
   input  wire  [16-1: 2] adc_dat_b_i        ,  // ADC CH2
   input  wire            adc_clk_p_i        ,  // ADC data clock
   input  wire            adc_clk_n_i        ,  // ADC data clock
   output wire  [ 2-1: 0] adc_clk_o          ,  // optional ADC clock source
   output wire            adc_cdcs_o         ,  // ADC clock duty cycle stabilizer
   // DAC
   output wire  [14-1: 0] dac_dat_o          ,  // DAC combined data
   output wire            dac_wrt_o          ,  // DAC write
   output wire            dac_sel_o          ,  // DAC channel select
   output wire            dac_clk_o          ,  // DAC clock
   output wire            dac_rst_o          ,  // DAC reset
   // PWM DAC
   output wire  [ 4-1: 0] dac_pwm_o          ,  // serial PWM DAC
   // XADC
   input  wire  [ 5-1: 0] vinp_i             ,  // voltages p
   input  wire  [ 5-1: 0] vinn_i             ,  // voltages n
   // Expansion connector
   inout  wire  [ 8-1: 0] exp_p_io           ,
   inout  wire  [ 8-1: 0] exp_n_io           ,
   // SATA connector
   output wire  [ 2-1: 0] daisy_p_o          ,  // line 1 is clock capable
   output wire  [ 2-1: 0] daisy_n_o          ,
   input  wire  [ 2-1: 0] daisy_p_i          ,  // line 1 is clock capable
   input  wire  [ 2-1: 0] daisy_n_i          ,
   // LED
   output wire  [ 8-1: 0] led_o       
);

//---------------------------------------------------------------------------------
//
//  Connections to PS

wire  [  4-1: 0] fclk               ; //[0]-125MHz, [1]-250MHz, [2]-50MHz, [3]-200MHz
wire  [  4-1: 0] frstn              ;

wire             ps_sys_clk         ;
wire             ps_sys_rstn        ;
wire  [ 32-1: 0] ps_sys_addr        ;
wire  [ 32-1: 0] ps_sys_wdata       ;
wire  [  4-1: 0] ps_sys_sel         ;
wire             ps_sys_wen         ;
wire             ps_sys_ren         ;
wire  [ 32-1: 0] ps_sys_rdata       ;
wire             ps_sys_err         ;
wire             ps_sys_ack         ;

// AXI masters
wire             axi1_clk    , axi0_clk    ;
wire             axi1_rstn   , axi0_rstn   ;
wire  [ 32-1: 0] axi1_waddr  , axi0_waddr  ;
wire  [ 64-1: 0] axi1_wdata  , axi0_wdata  ;
wire  [  8-1: 0] axi1_wsel   , axi0_wsel   ;
wire             axi1_wvalid , axi0_wvalid ;
wire  [  4-1: 0] axi1_wlen   , axi0_wlen   ;
wire             axi1_wfixed , axi0_wfixed ;
wire             axi1_werr   , axi0_werr   ;
wire             axi1_wrdy   , axi0_wrdy   ;

red_pitaya_ps i_ps (
  .FIXED_IO_mio       (  FIXED_IO_mio                ),
  .FIXED_IO_ps_clk    (  FIXED_IO_ps_clk             ),
  .FIXED_IO_ps_porb   (  FIXED_IO_ps_porb            ),
  .FIXED_IO_ps_srstb  (  FIXED_IO_ps_srstb           ),
  .FIXED_IO_ddr_vrn   (  FIXED_IO_ddr_vrn            ),
  .FIXED_IO_ddr_vrp   (  FIXED_IO_ddr_vrp            ),
  // DDR
  .DDR_addr      (DDR_addr    ),
  .DDR_ba        (DDR_ba      ),
  .DDR_cas_n     (DDR_cas_n   ),
  .DDR_ck_n      (DDR_ck_n    ),
  .DDR_ck_p      (DDR_ck_p    ),
  .DDR_cke       (DDR_cke     ),
  .DDR_cs_n      (DDR_cs_n    ),
  .DDR_dm        (DDR_dm      ),
  .DDR_dq        (DDR_dq      ),
  .DDR_dqs_n     (DDR_dqs_n   ),
  .DDR_dqs_p     (DDR_dqs_p   ),
  .DDR_odt       (DDR_odt     ),
  .DDR_ras_n     (DDR_ras_n   ),
  .DDR_reset_n   (DDR_reset_n ),
  .DDR_we_n      (DDR_we_n    ),

  .fclk_clk_o    (fclk        ),
  .fclk_rstn_o   (frstn       ),
  // ADC analog inputs
  .vinp_i        (vinp_i      ),  // voltages p
  .vinn_i        (vinn_i      ),  // voltages n
   // system read/write channel
  .sys_clk_o     (ps_sys_clk  ),  // system clock
  .sys_rstn_o    (ps_sys_rstn ),  // system reset - active low
  .sys_addr_o    (ps_sys_addr ),  // system read/write address
  .sys_wdata_o   (ps_sys_wdata),  // system write data
  .sys_sel_o     (ps_sys_sel  ),  // system write byte select
  .sys_wen_o     (ps_sys_wen  ),  // system write enable
  .sys_ren_o     (ps_sys_ren  ),  // system read enable
  .sys_rdata_i   (ps_sys_rdata),  // system read data
  .sys_err_i     (ps_sys_err  ),  // system error indicator
  .sys_ack_i     (ps_sys_ack  ),  // system acknowledge signal
  // AXI masters
  .axi1_clk_i    (axi1_clk    ),  .axi0_clk_i    (axi0_clk    ),  // global clock
  .axi1_rstn_i   (axi1_rstn   ),  .axi0_rstn_i   (axi0_rstn   ),  // global reset
  .axi1_waddr_i  (axi1_waddr  ),  .axi0_waddr_i  (axi0_waddr  ),  // system write address
  .axi1_wdata_i  (axi1_wdata  ),  .axi0_wdata_i  (axi0_wdata  ),  // system write data
  .axi1_wsel_i   (axi1_wsel   ),  .axi0_wsel_i   (axi0_wsel   ),  // system write byte select
  .axi1_wvalid_i (axi1_wvalid ),  .axi0_wvalid_i (axi0_wvalid ),  // system write data valid
  .axi1_wlen_i   (axi1_wlen   ),  .axi0_wlen_i   (axi0_wlen   ),  // system write burst length
  .axi1_wfixed_i (axi1_wfixed ),  .axi0_wfixed_i (axi0_wfixed ),  // system write burst type (fixed / incremental)
  .axi1_werr_o   (axi1_werr   ),  .axi0_werr_o   (axi0_werr   ),  // system write error
  .axi1_wrdy_o   (axi1_wrdy   ),  .axi0_wrdy_o   (axi0_wrdy   )   // system write ready
);

////////////////////////////////////////////////////////////////////////////////
// system bus decoder & multiplexer (it breaks memory addresses into 8 regions)
////////////////////////////////////////////////////////////////////////////////

wire              sys_clk   = ps_sys_clk  ;
wire              sys_rstn  = ps_sys_rstn ;
wire  [  32-1: 0] sys_addr  = ps_sys_addr ;
wire  [  32-1: 0] sys_wdata = ps_sys_wdata;
wire  [   4-1: 0] sys_sel   = ps_sys_sel  ;
wire  [8   -1: 0] sys_wen   ;
wire  [8   -1: 0] sys_ren   ;
wire  [8*32-1: 0] sys_rdata ;
wire  [8* 1-1: 0] sys_err   ;
wire  [8* 1-1: 0] sys_ack   ;
wire  [8   -1: 0] sys_cs    ;

assign sys_cs = 8'h01 << sys_addr[22:20];

assign sys_wen = sys_cs & {8{ps_sys_wen}};
assign sys_ren = sys_cs & {8{ps_sys_ren}};

assign ps_sys_rdata = sys_rdata[sys_addr[22:20]*32+:32];

assign ps_sys_err   = |(sys_cs & sys_err);
assign ps_sys_ack   = |(sys_cs & sys_ack);

// unused system bus slave ports

assign sys_rdata[5*32+:32] = 32'h0; 
assign sys_err  [5       ] =  1'b0;
assign sys_ack  [5       ] =  1'b1;

assign sys_rdata[6*32+:32] = 32'h0; 
assign sys_err  [6       ] =  1'b0;
assign sys_ack  [6       ] =  1'b1;

assign sys_rdata[7*32+:32] = 32'h0; 
assign sys_err  [7       ] =  1'b0;
assign sys_ack  [7       ] =  1'b1;

////////////////////////////////////////////////////////////////////////////////
// local signals
////////////////////////////////////////////////////////////////////////////////

// PLL signals
wire                  adc_clk_in;
wire                  pll_adc_clk;
wire                  pll_dac_clk_1x;
wire                  pll_dac_clk_2x;
wire                  pll_dac_clk_2p;
wire                  pll_clk_adc_2x;
wire                  pll_pwm_clk;
wire                  pll_locked;

// fast serial signals
wire                  ser_clk ;

// PWM clock and reset
wire                  pwm_clk ;
reg                   pwm_rstn;

// ADC signals
wire                  adc_clk, adc_clk_2x;
reg                   adc_rstn;
reg          [14-1:0] adc_dat_a, adc_dat_b;
wire  signed [14-1:0] adc_a    , adc_b    ;

// DAC signals
wire                  dac_clk_1x;
wire                  dac_clk_2x;
wire                  dac_clk_2p;
reg                   dac_rst;
reg          [14-1:0] dac_dat_a, dac_dat_b;
wire         [14-1:0] dac_a    , dac_b    ;
wire  signed [15-1:0] dac_a_sum, dac_b_sum;

// ASG
wire  signed [14-1:0] asg_a    , asg_b    ;

// PID
wire  signed [14-1:0] pid_a    , pid_b    ;

// configuration
wire                  digital_loop;

////////////////////////////////////////////////////////////////////////////////
// PLL (clock and reaset)
////////////////////////////////////////////////////////////////////////////////

// diferential clock input
IBUFDS i_clk (.I (adc_clk_p_i), .IB (adc_clk_n_i), .O (adc_clk_in));  // differential clock input

red_pitaya_pll pll (
  // inputs
  .clk         (adc_clk_in),  // clock
  .rstn        (frstn[0]  ),  // reset - active low
  // output clocks
  .clk_adc     (pll_adc_clk   ),  // ADC clock
  .clk_dac_1x  (pll_dac_clk_1x),  // DAC clock 125MHz
  .clk_dac_2x  (pll_dac_clk_2x),  // DAC clock 250MHz
  .clk_dac_2p  (pll_dac_clk_2p),  // DAC clock 250MHz -45DGR
  .clk_adc_2x  (pll_clk_adc_2x),  // fast serial clock
  .clk_pwm     (pll_pwm_clk   ),  // PWM clock
  // status outputs
  .pll_locked  (pll_locked)
);

BUFG bufg_adc_clk    (.O (adc_clk   ), .I (pll_adc_clk   ));
BUFG bufg_dac_clk_1x (.O (dac_clk_1x), .I (pll_dac_clk_1x));
BUFG bufg_dac_clk_2x (.O (dac_clk_2x), .I (pll_dac_clk_2x));
BUFG bufg_dac_clk_2p (.O (dac_clk_2p), .I (pll_dac_clk_2p));
BUFG bufg_ser_clk    (.O (adc_clk_2x), .I (pll_clk_adc_2x));
BUFG bufg_pwm_clk    (.O (pwm_clk   ), .I (pll_pwm_clk   ));

// ADC reset (active low) 
always @(posedge adc_clk)
adc_rstn <=  frstn[0] &  pll_locked;

// DAC reset (active high)
always @(posedge dac_clk_1x)
dac_rst  <= ~frstn[0] | ~pll_locked;

// PWM reset (active low)
always @(posedge pwm_clk)
pwm_rstn <=  frstn[0] &  pll_locked;

////////////////////////////////////////////////////////////////////////////////
// ADC IO
////////////////////////////////////////////////////////////////////////////////

// generating ADC clock is disabled
assign adc_clk_o = 2'b10;

// ADC clock duty cycle stabilizer is enabled
assign adc_cdcs_o = 1'b1 ;

// IO block registers should be used here
// lowest 2 bits reserved for 16bit ADC
always @(posedge adc_clk)
begin
  adc_dat_a <= adc_dat_a_i[16-1:2];
  adc_dat_b <= adc_dat_b_i[16-1:2];
end
    
// transform into 2's complement (negative slope)
assign adc_a = digital_loop ? dac_a : {adc_dat_a[14-1], ~adc_dat_a[14-2:0]};
assign adc_b = digital_loop ? dac_b : {adc_dat_b[14-1], ~adc_dat_b[14-2:0]};

////////////////////////////////////////////////////////////////////////////////
// DAC IO
////////////////////////////////////////////////////////////////////////////////

// // JD: Added a manual offset register for the dac outputs, at addresses 0x4050_0000 and 0x4050_0004:
// // manual output registers which add to the dac output value:


// output registers + signed to unsigned (also to negative slope)
always @(posedge dac_clk_1x)
begin
  dac_dat_a <= {dac_a[14-1], ~dac_a[14-2:0]};
  dac_dat_b <= {dac_b[14-1], ~dac_b[14-2:0]};
end

// DDR outputs
ODDR oddr_dac_clk          (.Q(dac_clk_o), .D1(1'b0     ), .D2(1'b1     ), .C(dac_clk_2p), .CE(1'b1), .R(1'b0   ), .S(1'b0));
ODDR oddr_dac_wrt          (.Q(dac_wrt_o), .D1(1'b0     ), .D2(1'b1     ), .C(dac_clk_2x), .CE(1'b1), .R(1'b0   ), .S(1'b0));
ODDR oddr_dac_sel          (.Q(dac_sel_o), .D1(1'b1     ), .D2(1'b0     ), .C(dac_clk_1x), .CE(1'b1), .R(dac_rst), .S(1'b0));
ODDR oddr_dac_rst          (.Q(dac_rst_o), .D1(dac_rst  ), .D2(dac_rst  ), .C(dac_clk_1x), .CE(1'b1), .R(1'b0   ), .S(1'b0));
ODDR oddr_dac_dat [14-1:0] (.Q(dac_dat_o), .D1(dac_dat_b), .D2(dac_dat_a), .C(dac_clk_1x), .CE(1'b1), .R(dac_rst), .S(1'b0));



//---------------------------------------------------------------------------------
//  Digital-PLL module (2 inputs, 2 outputs)
wire signed [15:0] ADCraw0, ADCraw1;
wire signed [15:0] DACout0, DACout1;
wire [16-1:0] LoggerData;
wire LoggerData_clk_enable;
wire LoggerIsWriting;

assign ADCraw0 = {adc_a, 2'b0};
assign ADCraw1 = {adc_b, 2'b0};
assign dac_a = DACout0[16-1:2];   // converts 16 bits DACout to 14 bits for dac_a
//assign dac_b = DACout1[16-1:2];   // converts 16 bits DACout to 14 bits for dac_b

wire dpll_rst = 1'b0; // I don't know if we can use the RedPitaya's reset because I don't know if it is clock-synchronous or not. In any case, it does not matter because we have the sys_bus driven resets.

dpll_wrapper dpll_wrapper_inst (
  
  .clk1                    (  adc_clk                    ), // global clock, designed for 100 MHz clock rate
  .clk1_timesN             (  adc_clk_2x                 ), // this should be N times the clock, phase-locked to clk1, N matching what was input in the FIR compiler for fir_compiler_minimumphase_N_times_clk
  .rst                     (  dpll_rst                   ), // currently only use the resets driven by the system bus

  // analog data input/output interface
  .ADCraw0                 (  ADCraw0                    ),
  .ADCraw1                 (  ADCraw1                    ),
  .DACout0                 (  DACout0                    ),
  .DACout1                 (  DACout1                    ),

  // Data logger port:
  .LoggerData              (  LoggerData                 ),
  .LoggerData_clk_enable   (  LoggerData_clk_enable      ),
  .LoggerIsWriting         (  LoggerIsWriting            ),

  // System bus
  .sys_addr                (  sys_addr                   ),  // address
  .sys_wdata               (  sys_wdata                  ),  // write data
  .sys_sel                 (  sys_sel                    ),  // write byte select
  .sys_wen                 (  sys_wen[0]                 ),  // write enable
  .sys_ren                 (  sys_ren[0]                 ),  // read enable
  .sys_rdata               (  sys_rdata[ 0*32+31: 0*32]  ),  // read data
  .sys_err                 (  sys_err[0]                 ),  // error indicator
  .sys_ack                 (  sys_ack[0]                 )   // acknowledge signal

);

// // ---------------------------------------------------------------------------------
// // For testing the N-times clk FIR filter:
// reg signed [16-1:0] fir_test_data;

// N_times_clk_FIR_wrapper N_times_clk_FIR_wrapper_inst (
//   // these two clocks need to be phase-locked to have a common edge (0 phase difference at the rising edges of clk_times_1)
//   .clk_times_1    (  adc_clk        ),
//   .clk_times_N    (  adc_clk_2x     ),
  
//   // these two signals are on the clk_times_1 clock domain
//   .data_in        (  fir_test_data  ),
//   .data_out       (  LoggerData     )

//   );
// assign LoggerData_clk_enable = 1'b1;

// always @(posedge adc_clk)
// begin
//   if (LoggerIsWriting) begin
//     fir_test_data <= 16'd1000;
//   end
//   else begin
//     fir_test_data <= 16'd0;
//   end
// end

//---------------------------------------------------------------------------------
// BRAM-based data logger, replaces the Red Pitaya oscilloscope application, but has much simpler behavior:
// The write port is directly controlled by the DPLL module, while the reads happen through the Zynq sys_bus

// // for testing independently of the DPLL module:
// assign LoggerData = adc_a;
// assign LoggerData_clk_enable = 1'b1;

ram_data_logger ram_data_logger_i (
  .clk                  (  adc_clk                    ),
  
  // data input interface
  .data_in              (  LoggerData                 ),
  .data_in_clk_enable   (  LoggerData_clk_enable      ),
  // control interface
  .is_writing           (  LoggerIsWriting            ),
  
  // CPU interface
  .sys_addr             (  sys_addr                   ),  // address
  .sys_wdata            (  sys_wdata                  ),  // write data
  .sys_sel              (  sys_sel                    ),  // write byte select
  .sys_wen              (  sys_wen[1]                 ),  // write enable
  .sys_ren              (  sys_ren[1]                 ),  // read enable
  .sys_rdata            (  sys_rdata[ 1*32+31: 1*32]  ),  // read data
  .sys_err              (  sys_err[1]                 ),  // error indicator
  .sys_ack              (  sys_ack[1]                 )   // acknowledge signal


  );


//---------------------------------------------------------------------------------
//  Internal VCO for testing purposes:
wire signed [16-1:0] vco_cosine_out;
wire signed [16-1:0] vco_sine_out;

reg  signed [48-1:0] vco_frequency;

always @(posedge adc_clk)
begin
  // gain was determined to mimick ~3e8 Hz/V of VCO gain, using:
  // log2(3e8/(125e6/2^48 * 2^15/1))
  // offset is equal to dec2bin(20e6/100e6 * 2^48, 48)
  vco_frequency <= ($signed(DACout0)<<<34) + $signed(48'b001100110011001100110011001100110011001100110011);
end

internal_vco internal_vco_i (

  .clk             (  adc_clk                    ),

  // frequency in counts: analog frequency is equal to: frequency/2^48*clock frequency (currently 125 MHz)
  .frequency       (  vco_frequency              ),

   // System bus, address starts at 0x4X20_0000
  .sys_addr        (  sys_addr                   ),  // address
  .sys_wdata       (  sys_wdata                  ),  // write data
  .sys_sel         (  sys_sel                    ),  // write byte select
  .sys_wen         (  sys_wen[2]                 ),  // write enable
  .sys_ren         (  sys_ren[2]                 ),  // read enable
  .sys_rdata       (  sys_rdata[ 2*32+31: 2*32]  ),  // read data
  .sys_err         (  sys_err[2]                 ),  // error indicator
  .sys_ack         (  sys_ack[2]                 ),  // acknowledge signal


  .cosine_out      (  vco_cosine_out             ),
  .sine_out        (  vco_sine_out               )

  );
assign dac_b = vco_cosine_out[16-1:2];

//---------------------------------------------------------------------------------
//  House Keeping

wire  [  8-1: 0] exp_p_in , exp_n_in ;
wire  [  8-1: 0] exp_p_out, exp_n_out;
wire  [  8-1: 0] exp_p_dir, exp_n_dir;

red_pitaya_hk i_hk (
  // system signals
  .clk_i           (  adc_clk                    ),  // clock
  .rstn_i          (  adc_rstn                   ),  // reset - active low
  // LED
  .led_o           (  led_o                      ),  // LED output
  // global configuration
  .digital_loop    (  digital_loop               ),
  // Expansion connector
  .exp_p_dat_i     (  exp_p_in                   ),  // input data
  .exp_p_dat_o     (  exp_p_out                  ),  // output data
  .exp_p_dir_o     (  exp_p_dir                  ),  // 1-output enable
  .exp_n_dat_i     (  exp_n_in                   ),
  .exp_n_dat_o     (  exp_n_out                  ),
  .exp_n_dir_o     (  exp_n_dir                  ),
   // System bus
  .sys_addr        (  sys_addr                   ),  // address
  .sys_wdata       (  sys_wdata                  ),  // write data
  .sys_sel         (  sys_sel                    ),  // write byte select
  .sys_wen         (  sys_wen[3]                 ),  // write enable
  .sys_ren         (  sys_ren[3]                 ),  // read enable
  .sys_rdata       (  sys_rdata[ 3*32+31: 3*32]  ),  // read data
  .sys_err         (  sys_err[3]                 ),  // error indicator
  .sys_ack         (  sys_ack[3]                 )   // acknowledge signal
);

IOBUF i_iobufp [8-1:0] (.O(exp_p_in), .IO(exp_p_io), .I(exp_p_out), .T(~exp_p_dir) );
IOBUF i_iobufn [8-1:0] (.O(exp_n_in), .IO(exp_n_io), .I(exp_n_out), .T(~exp_n_dir) );



// ---------------------------------------------------------------------------------
//  Oscilloscope application
// JDD: I kept this here just because it seems like we need to keep the axi0 and axi1 modules,
// otherwise the Zynq PS hangs up everytime we try to access the FPGA's address space.
// Eventually I should figure out how to properly remove them without this lock-up problem.
// It could simply be related to the fact that axi0_clk and axi1_clk are in fact connected to adc_clk inside this module,
// but it could also be that we need to 'ack' transactions in some manner which is implemented by the axi-fifos inside...

wire trig_asg_out ;

red_pitaya_scope i_scope (
  // ADC
  // .adc_a_i         (  adc_a                      ),  // CH 1
  // .adc_b_i         (  adc_b                      ),  // CH 2
  .adc_clk_i       (  adc_clk                    ),  // clock
  .adc_rstn_i      (  adc_rstn                   ),  // reset - active low
  // .trig_ext_i      (  exp_p_in[0]                ),  // external trigger
  // .trig_asg_i      (  trig_asg_out               ),  // ASG trigger
  // AXI0 master                 // AXI1 master
  .axi0_clk_o    (axi0_clk   ),  .axi1_clk_o    (axi1_clk   ),
  .axi0_rstn_o   (axi0_rstn  ),  .axi1_rstn_o   (axi1_rstn  ),
  .axi0_waddr_o  (axi0_waddr ),  .axi1_waddr_o  (axi1_waddr ),
  .axi0_wdata_o  (axi0_wdata ),  .axi1_wdata_o  (axi1_wdata ),
  .axi0_wsel_o   (axi0_wsel  ),  .axi1_wsel_o   (axi1_wsel  ),
  .axi0_wvalid_o (axi0_wvalid),  .axi1_wvalid_o (axi1_wvalid),
  .axi0_wlen_o   (axi0_wlen  ),  .axi1_wlen_o   (axi1_wlen  ),
  .axi0_wfixed_o (axi0_wfixed),  .axi1_wfixed_o (axi1_wfixed),
  .axi0_werr_i   (axi0_werr  ),  .axi1_werr_i   (axi1_werr  ),
  .axi0_wrdy_i   (axi0_wrdy  ),  .axi1_wrdy_i   (axi1_wrdy  )
  // // System bus
  // .sys_addr        (  sys_addr                   ),  // address
  // .sys_wdata       (  sys_wdata                  ),  // write data
  // .sys_sel         (  sys_sel                    ),  // write byte select
  // .sys_wen         (  sys_wen[1]                 ),  // write enable
  // .sys_ren         (  sys_ren[1]                 ),  // read enable
  // .sys_rdata       (  sys_rdata[ 1*32+31: 1*32]  ),  // read data
  // .sys_err         (  sys_err[1]                 ),  // error indicator
  // .sys_ack         (  sys_ack[1]                 )   // acknowledge signal
);



//---------------------------------------------------------------------------------
//  Daisy chain
//  simple communication module

assign daisy_p_o = 1'bz;
assign daisy_n_o = 1'bz;

endmodule

